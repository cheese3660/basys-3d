library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package basys3d_arithmetic is
    type divider_array_t is array(natural range <>) of signed; 
end basys3d_arithmetic;